library ieee;
use ieee.std_logic_1164.all;

package fsm_package is
    type state_type is (S01, S11, S10, S00);
end package;