library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package fsm_package is
    type state_type is (S0, S1, S2);
end package;

package body fsm_package is
end package body;